module Perm(
	input [4:0] perm_in_5,
	input [8:0] perm_in_9,
	output [4:0] perm_out
	);
	
	wire [4:0] ind_perm_out;
	
	always @(*) begin
			
	end
endmodule
