module perm_stage(

	);

endmodule